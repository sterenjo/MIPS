-- Ifetch module (provides the PC and instruction 
--memory for the MIPS computer)
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY Ifetch IS
	PORT(	SIGNAL Instruction 		: OUT	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        	SIGNAL PC_plus_4_out 	: OUT	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
        	SIGNAL Add_result 		: IN 	STD_LOGIC_VECTOR( 7 DOWNTO 0 );
        	SIGNAL beq,bne 			: IN 	STD_LOGIC;
        	SIGNAL Zero 			: IN 	STD_LOGIC;
      		SIGNAL PC_out 			: OUT	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
        	SIGNAL clock			: IN 	STD_LOGIC;
			SIGNAL reset 			: IN 	STD_LOGIC;
			SIGNAL J			 	: IN 	STD_LOGIC;
			SIGNAL JR			 	: IN 	STD_LOGIC;
			SIGNAL read_data_1 		: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 ));
END Ifetch;

ARCHITECTURE behavior OF Ifetch IS
	SIGNAL PC, PC_plus_4 	 : STD_LOGIC_VECTOR( 9 DOWNTO 0 );
	SIGNAL next_PC, Mem_Addr : STD_LOGIC_VECTOR( 7 DOWNTO 0 );
	SIGNAL modelsim : boolean;
	
BEGIN 
						--ROM for Instruction Memory
inst_memory: altsyncram
modelsim <= TRUE;
	
	GENERIC MAP (
		operation_mode => "ROM",
		width_a => 32,
		widthad_a => 8,
		lpm_type => "altsyncram",
		outdata_reg_a => "UNREGISTERED",
		init_file => "C:\TestPrograms\ModelSim\L1_Cache\asm_ver1\program.hex",
		intended_device_family => "Cyclone"
	)
	PORT MAP (
		clock0     => clock,
		address_a 	=> Mem_Addr, 
		q_a 			=> Instruction );
		
		
					-- Instructions always start on word address - not byte
		PC(1 DOWNTO 0) <= "00";
		
					-- copy output signals - allows read inside module
		PC_out 			<= PC;
		PC_plus_4_out 	<= PC_plus_4;
		
						-- send address to inst. memory address registerIF
		if (modelsim = TRUE) generate
			Mem_Addr <= Next_PC;
		end generate;
		
		if (modelsim = FALSE ) generate
			Mem_Addr <= Next_PC & "00";
		end generate;
		
						-- Adder to increment PC by 4        
      	PC_plus_4( 9 DOWNTO 2 )  <= PC( 9 DOWNTO 2 ) + 1;
       	PC_plus_4( 1 DOWNTO 0 )  <= "00";
		
						-- Mux to select Branch Address or PC + 4        
		Next_PC  <= X"00" WHEN Reset = '1' 
			ELSE    Add_result WHEN ( ( ( beq = '1' ) AND ( Zero = '1' ) ) OR ( ( bne = '1' ) AND ( Zero = '0' ) )) -- Branch (jump = '1'?)
			ELSE  	Instruction(7 DOWNTO 0) WHEN J = '1' 	 --- J instuction ---
			ELSE 	read_data_1(9 DOWNTO 2) WHEN JR = '1'  --- JR instuction ---
			ELSE    PC_plus_4  ( 9 DOWNTO 2 );
			
	PROCESS
		BEGIN
			WAIT UNTIL ( clock'EVENT ) AND ( clock = '1' );
			IF reset = '1' THEN
				   PC( 9 DOWNTO 2) <= "00000000" ; 
			ELSE 
				   PC( 9 DOWNTO 2 ) <= next_PC;
			END IF;
	END PROCESS;
END behavior;


